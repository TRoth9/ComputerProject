module Accumulator	(output reg [7:0] Acc_out,
							 input [7:0] Bus_in,
							 input OE,
							 input WE,
							 input CLK,
							 input RESET);
		
		reg [7:0] Acc;
		
		always @(Acc_out or OE or WE) begin
			if (!OE) begin
				Acc_out <= 8b'00000000;
			end
		end
		
		always @(posedge CLK or posedge RESET) begin
				if (RESET) begin
					Acc <= 8b'00000000;
					Acc_out <= 8b'00000000;
				end					
				else if (WE) begin
					Acc <= Bus_in;
				end
				else if (OE) begin
					Acc_out <= Acc;
				end
		end

endmodule